// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
`ifndef CL_NOVA_DEFINES
`define CL_NOVA_DEFINES
//Put module name of the CL design here.  This is used to instantiate in top.sv
`define CL_NAME cl_top

//Highly recommeneded.  For lib FIFO block, uses less async reset (take advantage of
// FPGA flop init capability).  This will help with routing resources.
`define FPGA_LESS_RST

// Uncomment to disable Virtual JTAG
`define DISABLE_VJTAG_DEBUG

//Must have this define or will get syntax errors.  Curretly XDMA not supported.
// `define NO_XDMA
`endif 
